x"20", x"00", x"68", x"8e", x"20", x"40", x"48", x"02", x"20", x"00", x"68", x"ae", 